CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
1093 99 1909 1007
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
1261 195 1374 292
9437202 0
0
6 Title:
5 Name:
0
0
0
29
13 Logic Switch~
5 109 485 0 1 11
0 27
0
0 0 21360 0
2 0V
-6 -16 8 -8
6 Enable
-20 -26 22 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 512 0 0 -1 0
1 V
5130 0 0
2
43535.1 0
0
13 Logic Switch~
5 109 439 0 1 11
0 10
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 D8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
391 0 0
2
43535.1 0
0
13 Logic Switch~
5 108 265 0 1 11
0 22
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 D4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3124 0 0
2
43535.1 3
0
13 Logic Switch~
5 108 300 0 1 11
0 21
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 D5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3421 0 0
2
43535.1 2
0
13 Logic Switch~
5 110 353 0 1 11
0 20
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 D6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8157 0 0
2
43535.1 1
0
13 Logic Switch~
5 110 388 0 1 11
0 19
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 D7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5572 0 0
2
43535.1 0
0
13 Logic Switch~
5 107 177 0 1 11
0 24
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 D2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8901 0 0
2
43535.1 1
0
13 Logic Switch~
5 107 212 0 1 11
0 23
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 D3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7361 0 0
2
43535.1 0
0
13 Logic Switch~
5 105 124 0 1 11
0 25
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 D1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4747 0 0
2
43535.1 0
0
13 Logic Switch~
5 105 89 0 1 11
0 26
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 D0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
972 0 0
2
43535.1 0
0
5 4049~
219 158 262 0 2 22
0 22 15
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U6B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 6 0
1 U
3472 0 0
2
43535.1 3
0
5 4049~
219 157 296 0 2 22
0 21 16
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U6A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 6 0
1 U
9998 0 0
2
43535.1 2
0
5 4049~
219 157 386 0 2 22
0 19 17
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U5F
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 5 0
1 U
3536 0 0
2
43535.1 1
0
5 4049~
219 158 352 0 2 22
0 20 18
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U5E
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 5 0
1 U
4597 0 0
2
43535.1 0
0
5 4049~
219 153 177 0 2 22
0 24 13
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U5D
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 5 0
1 U
3835 0 0
2
43535.1 1
0
5 4049~
219 152 211 0 2 22
0 23 14
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U5C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 5 0
1 U
3670 0 0
2
43535.1 0
0
5 4049~
219 152 121 0 2 22
0 25 12
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U5B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 5 0
1 U
5616 0 0
2
43535.1 0
0
5 4049~
219 153 87 0 2 22
0 26 11
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U5A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 5 0
1 U
9323 0 0
2
43535.1 0
0
9 2-In AND~
219 660 257 0 3 22
0 28 2 29
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4B
-12 -25 9 -17
11 Even Output
-40 -45 37 -37
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 2 4 0
1 U
317 0 0
2
43535.1 0
0
6 74266~
219 538 266 0 3 22
0 9 10 2
0
0 0 624 0
7 74LS266
-24 -24 25 -16
3 U3A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3108 0 0
2
43535.1 0
0
9 2-In AND~
219 659 124 0 3 22
0 30 31 32
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4A
-12 -25 9 -17
11 Even Output
-40 -45 37 -37
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 1 4 0
1 U
4299 0 0
2
43535.1 0
0
6 74136~
219 539 134 0 3 22
0 10 9 33
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U2D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 4 2 0
1 U
9672 0 0
2
43535.1 0
0
6 74136~
219 437 219 0 3 22
0 8 7 9
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U2C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
7876 0 0
2
43535.1 0
0
6 74136~
219 218 363 0 3 22
0 18 17 5
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U2B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
6369 0 0
2
43535.1 2
0
6 74136~
219 326 310 0 3 22
0 6 5 7
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U2A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
9172 0 0
2
43535.1 1
0
6 74136~
219 218 274 0 3 22
0 15 16 6
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U1D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
7100 0 0
2
43535.1 0
0
6 74136~
219 324 137 0 3 22
0 3 4 8
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U1C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
3820 0 0
2
43535.1 0
0
6 74136~
219 216 190 0 3 22
0 13 14 4
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U1B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
7678 0 0
2
43535.1 0
0
6 74136~
219 216 101 0 3 22
0 11 12 3
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U1A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
961 0 0
2
43535.1 0
0
30
1 0 0 0 0 16 0 19 0 0 3 2
636 248
622 248
2 3 0 0 0 0 0 21 22 0 0 4
635 133
580 133
580 134
572 134
1 1 0 0 0 0 0 1 21 0 0 4
121 485
622 485
622 115
635 115
3 2 2 0 0 4224 0 20 19 0 0 2
577 266
636 266
1 3 3 0 0 4224 0 27 29 0 0 4
308 128
257 128
257 101
249 101
2 3 4 0 0 4224 0 27 28 0 0 4
308 146
257 146
257 190
249 190
2 3 5 0 0 4224 0 25 24 0 0 4
310 319
259 319
259 363
251 363
1 3 6 0 0 4224 0 25 26 0 0 4
310 301
259 301
259 274
251 274
2 3 7 0 0 8320 0 23 25 0 0 4
421 228
367 228
367 310
359 310
1 3 8 0 0 8320 0 23 27 0 0 4
421 210
365 210
365 137
357 137
1 0 9 0 0 8192 0 20 0 0 12 3
522 257
515 257
515 219
3 2 9 0 0 8320 0 23 22 0 0 4
470 219
515 219
515 143
523 143
2 0 10 0 0 4096 0 20 0 0 14 2
522 275
497 275
1 1 10 0 0 4224 0 2 22 0 0 4
121 439
497 439
497 125
523 125
2 1 11 0 0 4224 0 18 29 0 0 4
174 87
192 87
192 92
200 92
2 2 12 0 0 4224 0 17 29 0 0 4
173 121
192 121
192 110
200 110
2 1 13 0 0 4224 0 15 28 0 0 4
174 177
192 177
192 181
200 181
2 2 14 0 0 4224 0 16 28 0 0 4
173 211
192 211
192 199
200 199
2 1 15 0 0 4224 0 11 26 0 0 4
179 262
194 262
194 265
202 265
2 2 16 0 0 4224 0 12 26 0 0 4
178 296
194 296
194 283
202 283
2 2 17 0 0 4224 0 13 24 0 0 4
178 386
194 386
194 372
202 372
2 1 18 0 0 4224 0 14 24 0 0 4
179 352
194 352
194 354
202 354
1 1 19 0 0 4224 0 6 13 0 0 4
122 388
134 388
134 386
142 386
1 1 20 0 0 4224 0 5 14 0 0 4
122 353
135 353
135 352
143 352
1 1 21 0 0 4224 0 4 12 0 0 4
120 300
134 300
134 296
142 296
1 1 22 0 0 4224 0 3 11 0 0 4
120 265
135 265
135 262
143 262
1 1 23 0 0 4224 0 8 16 0 0 4
119 212
129 212
129 211
137 211
1 1 24 0 0 4224 0 7 15 0 0 2
119 177
138 177
1 1 25 0 0 4224 0 9 17 0 0 4
117 124
129 124
129 121
137 121
1 1 26 0 0 4224 0 10 18 0 0 4
117 89
130 89
130 87
138 87
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
