CircuitMaker Text
5.6
Probes: 1
L1_1
DC Sweep
0 534 355 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
150 100 30 150 10
1093 99 1909 1007
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
1261 195 2077 649
9961490 0
0
6 Title:
5 Name:
0
0
0
11
13 Logic Switch~
5 231 477 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7876 0 0
2
5.89884e-315 0
0
13 Logic Switch~
5 230 397 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6369 0 0
2
5.89884e-315 0
0
9 P-MESFET~
219 488 270 0 3 7
0 4 5 3
0
0 0 848 0
7 PMESFET
11 0 60 8
2 Q7
29 -10 43 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
122 0 0 0 0 0 0 0
1 Q
9172 0 0
2
43535.1 0
0
9 N-MESFET~
219 488 400 0 3 7
0 3 5 2
0
0 0 848 0
7 NMESFET
11 0 60 8
2 Q5
29 -10 43 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
90 0 0 0 0 0 0 0
1 Q
7100 0 0
2
43535.1 0
0
7 Ground~
168 350 523 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3820 0 0
2
5.89884e-315 0
0
2 +V
167 348 178 0 1 3
0 4
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7678 0 0
2
5.89884e-315 0
0
14 Logic Display~
6 579 332 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
961 0 0
2
5.89884e-315 0
0
9 N-MESFET~
219 342 477 0 3 7
0 8 6 2
0
0 0 848 0
7 NMESFET
11 0 60 8
2 Q4
29 -10 43 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
90 0 0 0 1 0 0 0
1 Q
3178 0 0
2
5.89884e-315 0
0
9 N-MESFET~
219 342 397 0 3 7
0 5 7 8
0
0 0 848 0
7 NMESFET
9 0 58 8
2 Q3
29 -10 43 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
90 0 0 0 1 0 0 0
1 Q
3409 0 0
2
5.89884e-315 0
0
9 P-MESFET~
219 430 264 0 3 7
0 4 6 5
0
0 0 848 512
7 PMESFET
-67 0 -18 8
2 Q2
-49 -10 -35 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
122 0 0 0 1 0 0 0
1 Q
3951 0 0
2
5.89884e-315 0
0
9 P-MESFET~
219 282 264 0 3 7
0 4 7 5
0
0 0 848 0
7 PMESFET
11 0 60 8
2 Q1
29 -10 43 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
122 0 0 0 1 0 0 0
1 Q
8885 0 0
2
5.89884e-315 0
0
16
1 0 3 0 0 8192 0 7 0 0 2 3
579 350
579 354
496 354
3 1 3 0 0 4240 0 3 4 0 0 2
496 288
496 382
1 0 4 0 0 8320 0 3 0 0 8 3
496 252
496 201
348 201
2 0 5 0 0 8192 0 4 0 0 5 3
475 400
467 400
467 337
0 2 5 0 0 4096 0 0 3 13 0 4
350 337
467 337
467 270
475 270
0 3 2 0 0 4224 0 0 4 7 0 3
350 509
496 509
496 418
1 3 2 0 0 128 0 5 8 0 0 2
350 517
350 495
1 0 4 0 0 0 0 6 0 0 14 2
348 187
348 238
0 2 6 0 0 12416 0 0 10 10 0 5
268 477
268 563
445 563
445 264
437 264
1 2 6 0 0 0 0 1 8 0 0 2
243 477
329 477
0 2 7 0 0 4224 0 0 11 12 0 3
261 397
261 264
269 264
1 2 7 0 0 0 0 2 9 0 0 2
242 397
329 397
1 0 5 0 0 0 0 9 0 0 15 2
350 379
350 290
1 1 4 0 0 128 0 11 10 0 0 4
290 246
290 238
416 238
416 246
3 3 5 0 0 8320 0 11 10 0 0 4
290 282
290 290
416 290
416 282
1 3 8 0 0 4224 0 8 9 0 0 2
350 459
350 415
0
0
2071 0 1
2 V3
0
2 V3
0 5 0.001
0
0 0 0
3 0 1 4
0 5e-06 2e-08 2e-08
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
