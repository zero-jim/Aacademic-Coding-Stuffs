CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
50 20 30 200 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
9
13 Logic Switch~
5 121 239 0 1 11
0 7
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
43283 0
0
13 Logic Switch~
5 128 168 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
391 0 0
2
43283 0
0
13 Logic Switch~
5 129 135 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3124 0 0
2
43283 0
0
13 Logic Switch~
5 130 99 0 1 11
0 9
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3421 0 0
2
43283 0
0
13 Logic Switch~
5 130 63 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
8157 0 0
2
43283 0
0
14 Logic Display~
6 449 191 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5572 0 0
2
43283 0
0
5 4049~
219 189 183 0 2 22
0 4 5
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U2B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 1 0
1 U
8901 0 0
2
43283 0
0
5 4049~
219 180 221 0 2 22
0 7 6
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U2A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 1 0
1 U
7361 0 0
2
43283 0
0
6 CD4512
77 294 173 0 14 29
0 4 7 7 5 5 7 6 6 2
9 8 7 7 3
0
0 0 4848 0
4 4512
-14 -60 14 -52
2 U1
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
146 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 9 7 6 5 4 3 2 1 13
12 11 15 10 14 9 7 6 5 4
3 2 1 13 12 11 15 10 14 0
65 0 0 0 0 0 0 0
1 U
4747 0 0
2
43283 0
0
17
0 9 2 0 0 8192 0 0 9 17 0 3
340 144
340 146
326 146
14 1 3 0 0 4224 0 9 6 0 0 2
326 209
449 209
0 1 4 0 0 8320 0 0 9 6 0 3
166 168
166 146
262 146
0 4 5 0 0 8192 0 0 9 5 0 3
213 182
213 173
262 173
2 5 5 0 0 8320 0 7 9 0 0 3
210 183
210 182
262 182
1 1 4 0 0 0 0 2 7 0 0 4
140 168
166 168
166 183
174 183
0 7 6 0 0 8192 0 0 9 8 0 3
237 210
237 200
262 200
2 8 6 0 0 4240 0 8 9 0 0 4
201 221
237 221
237 209
262 209
0 1 7 0 0 4096 0 0 8 14 0 3
152 239
152 221
165 221
0 2 7 0 0 0 0 0 9 11 0 3
254 165
254 155
262 155
0 3 7 0 0 4096 0 0 9 14 0 3
254 193
254 164
262 164
13 0 7 0 0 0 0 9 0 0 13 2
332 191
340 191
0 12 7 0 0 8192 0 0 9 14 0 5
254 239
254 224
340 224
340 182
332 182
1 6 7 0 0 4224 0 1 9 0 0 4
133 239
254 239
254 191
262 191
11 1 8 0 0 20608 0 9 5 0 0 6
326 164
350 164
350 146
350 146
350 63
142 63
10 1 9 0 0 12416 0 9 4 0 0 4
326 155
345 155
345 99
142 99
0 1 2 0 0 8320 0 0 3 0 0 4
340 164
340 117
141 117
141 135
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
