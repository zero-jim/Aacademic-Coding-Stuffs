CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
60 0 30 150 10
1093 99 1909 1007
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
1261 195 1374 292
9437202 0
0
6 Title:
5 Name:
0
0
0
12
13 Logic Switch~
5 130 179 0 1 11
0 2
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
43535.1 0
0
13 Logic Switch~
5 130 102 0 1 11
0 3
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
391 0 0
2
43535.1 0
0
5 4049~
219 211 179 0 2 22
0 2 8
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U2B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 512 6 2 2 0
1 U
3124 0 0
2
43535.1 0
0
5 4049~
219 212 101 0 2 22
0 3 9
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U2A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 512 6 1 2 0
1 U
3421 0 0
2
43535.1 0
0
9 2-In AND~
219 456 268 0 3 22
0 10 11 4
0
0 0 624 0
6 74LS08
-21 -24 21 -16
2 D3
-9 -25 5 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 4 1 0
1 U
8157 0 0
2
43535.1 1
0
9 2-In AND~
219 455 214 0 3 22
0 12 13 5
0
0 0 624 0
6 74LS08
-21 -24 21 -16
2 D2
-9 -25 5 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 3 1 0
1 U
5572 0 0
2
43535.1 0
0
9 2-In AND~
219 452 164 0 3 22
0 14 15 6
0
0 0 624 0
6 74LS08
-21 -24 21 -16
2 D1
-9 -25 5 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 2 1 0
1 U
8901 0 0
2
43535.1 0
0
9 2-In AND~
219 452 109 0 3 22
0 16 17 7
0
0 0 624 0
6 74LS08
-21 -24 21 -16
2 D0
-9 -25 5 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 1 1 0
1 U
7361 0 0
2
43535.1 0
0
14 Logic Display~
6 509 255 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4747 0 0
2
43535.1 0
0
14 Logic Display~
6 507 195 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
972 0 0
2
43535.1 0
0
14 Logic Display~
6 507 146 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3472 0 0
2
43535.1 0
0
14 Logic Display~
6 506 95 0 1 2
10 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9998 0 0
2
43535.1 0
0
14
1 0 0 0 0 0 0 6 0 0 2 2
431 205
191 205
0 1 0 0 0 0 0 0 5 9 0 3
191 179
191 259
432 259
1 0 0 0 0 16 0 7 0 0 4 4
428 155
189 155
189 156
174 156
0 2 0 0 0 0 0 0 5 10 0 3
174 102
174 277
432 277
2 0 0 0 0 0 0 7 0 0 6 2
428 173
420 173
2 2 0 0 0 0 0 3 8 0 0 4
232 179
420 179
420 118
428 118
1 0 0 0 0 0 0 8 0 0 8 3
428 100
409 100
409 101
2 2 0 0 0 0 0 4 6 0 0 4
233 101
410 101
410 223
431 223
1 1 2 0 0 4224 0 1 3 0 0 2
142 179
196 179
1 1 3 0 0 4224 0 2 4 0 0 4
142 102
188 102
188 101
197 101
3 1 4 0 0 4224 0 5 9 0 0 5
477 268
497 268
497 281
509 281
509 273
3 1 5 0 0 4224 0 6 10 0 0 5
476 214
495 214
495 221
507 221
507 213
3 1 6 0 0 4224 0 7 11 0 0 5
473 164
495 164
495 172
507 172
507 164
3 1 7 0 0 4224 0 8 12 0 0 5
473 109
494 109
494 121
506 121
506 113
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
