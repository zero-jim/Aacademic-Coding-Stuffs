CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 120 10
1093 99 1909 1007
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
1261 195 1374 292
9437202 0
0
6 Title:
5 Name:
0
0
0
37
5 4071~
219 415 871 0 3 22
0 5 4 2
0
0 0 608 0
4 4071
-7 -24 21 -16
3 U1D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 1 0
1 U
5130 0 0
2
43535.1 9
0
5 4030~
219 262 787 0 3 22
0 9 8 7
0
0 0 608 0
4 4030
-7 -24 21 -16
3 U4D
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 4 0
1 U
391 0 0
2
43535.1 8
0
5 4030~
219 348 795 0 3 22
0 7 6 3
0
0 0 608 0
4 4030
-7 -24 21 -16
3 U4C
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 4 0
1 U
3124 0 0
2
43535.1 7
0
5 4081~
219 359 894 0 3 22
0 9 8 4
0
0 0 608 0
4 4081
-7 -24 21 -16
3 U5D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 5 0
1 U
3421 0 0
2
43535.1 6
0
5 4081~
219 358 848 0 3 22
0 7 6 5
0
0 0 608 0
4 4081
-7 -24 21 -16
3 U5C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 5 0
1 U
8157 0 0
2
43535.1 5
0
14 Logic Display~
6 508 777 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5572 0 0
2
43535.1 4
0
14 Logic Display~
6 495 853 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8901 0 0
2
43535.1 3
0
13 Logic Switch~
5 168 778 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 A3
-8 -33 6 -25
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7361 0 0
2
43535.1 2
0
13 Logic Switch~
5 170 812 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 B3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4747 0 0
2
43535.1 1
0
13 Logic Switch~
5 167 612 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 B2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
972 0 0
2
43535.1 8
0
13 Logic Switch~
5 165 578 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 A2
-8 -33 6 -25
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3472 0 0
2
43535.1 7
0
14 Logic Display~
6 492 653 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9998 0 0
2
43535.1 6
0
14 Logic Display~
6 505 577 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3536 0 0
2
43535.1 5
0
5 4081~
219 355 648 0 3 22
0 7 6 5
0
0 0 608 0
4 4081
-7 -24 21 -16
3 U5B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 5 0
1 U
4597 0 0
2
43535.1 4
0
5 4081~
219 356 694 0 3 22
0 9 8 4
0
0 0 608 0
4 4081
-7 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 5 0
1 U
3835 0 0
2
43535.1 3
0
5 4030~
219 345 595 0 3 22
0 7 6 3
0
0 0 608 0
4 4030
-7 -24 21 -16
3 U4B
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 4 0
1 U
3670 0 0
2
43535.1 2
0
5 4030~
219 259 587 0 3 22
0 9 8 7
0
0 0 608 0
4 4030
-7 -24 21 -16
3 U4A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 4 0
1 U
5616 0 0
2
43535.1 1
0
5 4071~
219 412 671 0 3 22
0 5 4 2
0
0 0 608 0
4 4071
-7 -24 21 -16
3 U1C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 1 0
1 U
9323 0 0
2
43535.1 0
0
5 4071~
219 407 475 0 3 22
0 5 4 2
0
0 0 608 0
4 4071
-7 -24 21 -16
3 U1B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 1 0
1 U
317 0 0
2
43535.1 9
0
5 4030~
219 254 391 0 3 22
0 9 8 7
0
0 0 608 0
4 4030
-7 -24 21 -16
3 U2D
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 2 0
1 U
3108 0 0
2
43535.1 8
0
5 4030~
219 340 399 0 3 22
0 7 6 3
0
0 0 608 0
4 4030
-7 -24 21 -16
3 U2C
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 2 0
1 U
4299 0 0
2
43535.1 7
0
5 4081~
219 351 498 0 3 22
0 9 8 4
0
0 0 608 0
4 4081
-7 -24 21 -16
3 U3D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 3 0
1 U
9672 0 0
2
43535.1 6
0
5 4081~
219 350 452 0 3 22
0 7 6 5
0
0 0 608 0
4 4081
-7 -24 21 -16
3 U3C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 3 0
1 U
7876 0 0
2
43535.1 5
0
14 Logic Display~
6 500 381 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6369 0 0
2
43535.1 4
0
14 Logic Display~
6 487 457 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9172 0 0
2
43535.1 3
0
13 Logic Switch~
5 160 382 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 A1
-8 -33 6 -25
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7100 0 0
2
43535.1 2
0
13 Logic Switch~
5 162 416 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 B1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3820 0 0
2
43535.1 1
0
13 Logic Switch~
5 161 324 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
3 Cin
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7678 0 0
2
43535.1 0
0
13 Logic Switch~
5 162 217 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 B0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
961 0 0
2
43535.1 1
0
13 Logic Switch~
5 160 183 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 A0
-8 -33 6 -25
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3178 0 0
2
43535.1 2
0
14 Logic Display~
6 487 258 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3409 0 0
2
43535.1 3
0
14 Logic Display~
6 500 182 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3951 0 0
2
43535.1 4
0
5 4081~
219 350 253 0 3 22
0 7 6 5
0
0 0 608 0
4 4081
-7 -24 21 -16
3 U3B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 3 0
1 U
8885 0 0
2
43535.1 5
0
5 4081~
219 351 299 0 3 22
0 9 8 4
0
0 0 608 0
4 4081
-7 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 3 0
1 U
3780 0 0
2
43535.1 6
0
5 4030~
219 340 200 0 3 22
0 7 6 3
0
0 0 608 0
4 4030
-7 -24 21 -16
3 U2B
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 2 0
1 U
9265 0 0
2
43535.1 7
0
5 4030~
219 254 192 0 3 22
0 9 8 7
0
0 0 608 0
4 4030
-7 -24 21 -16
3 U2A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 2 0
1 U
9442 0 0
2
43535.1 8
0
5 4071~
219 407 276 0 3 22
0 5 4 2
0
0 0 608 0
4 4071
-7 -24 21 -16
3 U1A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 1 0
1 U
9424 0 0
2
43535.1 9
0
48
3 1 2 0 0 0 0 1 7 0 0 2
448 871
495 871
3 1 3 0 0 0 0 3 6 0 0 2
381 795
508 795
3 2 4 0 0 0 0 4 1 0 0 3
380 894
380 880
402 880
3 1 5 0 0 0 0 5 1 0 0 4
379 848
380 848
380 862
402 862
0 2 6 0 0 0 0 0 5 7 0 3
304 804
304 857
334 857
0 1 7 0 0 0 0 0 5 8 0 3
297 788
297 839
334 839
0 2 6 0 0 16 0 0 3 13 0 5
460 671
460 755
304 755
304 804
332 804
3 1 7 0 0 0 0 2 3 0 0 5
295 787
295 788
297 788
297 786
332 786
0 2 8 0 0 0 0 0 4 11 0 3
199 812
199 903
335 903
0 1 9 0 0 0 0 0 4 12 0 3
216 778
216 885
335 885
1 2 8 0 0 0 0 9 2 0 0 4
182 812
224 812
224 796
246 796
1 1 9 0 0 0 0 8 2 0 0 2
180 778
246 778
3 1 2 0 0 0 0 18 12 0 0 2
445 671
492 671
3 1 3 0 0 0 0 16 13 0 0 2
378 595
505 595
3 2 4 0 0 0 0 15 18 0 0 3
377 694
377 680
399 680
3 1 5 0 0 0 0 14 18 0 0 4
376 648
377 648
377 662
399 662
0 2 6 0 0 0 0 0 14 19 0 3
301 604
301 657
331 657
0 1 7 0 0 0 0 0 14 20 0 3
294 588
294 639
331 639
0 2 6 0 0 0 0 0 16 25 0 5
451 475
451 552
301 552
301 604
329 604
3 1 7 0 0 0 0 17 16 0 0 5
292 587
292 588
294 588
294 586
329 586
0 2 8 0 0 0 0 0 15 23 0 3
196 612
196 703
332 703
0 1 9 0 0 0 0 0 15 24 0 3
213 578
213 685
332 685
1 2 8 0 0 0 0 10 17 0 0 4
179 612
221 612
221 596
243 596
1 1 9 0 0 0 0 11 17 0 0 2
177 578
243 578
3 1 2 0 0 0 0 19 25 0 0 2
440 475
487 475
3 1 3 0 0 0 0 21 24 0 0 2
373 399
500 399
3 2 4 0 0 0 0 22 19 0 0 3
372 498
372 484
394 484
3 1 5 0 0 0 0 23 19 0 0 4
371 452
372 452
372 466
394 466
0 2 6 0 0 0 0 0 23 31 0 3
296 408
296 461
326 461
0 1 7 0 0 0 0 0 23 32 0 3
289 392
289 443
326 443
0 2 6 0 0 0 0 0 21 37 0 5
462 276
462 358
295 358
295 408
324 408
3 1 7 0 0 0 0 20 21 0 0 5
287 391
287 392
289 392
289 390
324 390
0 2 8 0 0 0 0 0 22 35 0 3
191 416
191 507
327 507
0 1 9 0 0 0 0 0 22 36 0 3
208 382
208 489
327 489
1 2 8 0 0 0 0 27 20 0 0 4
174 416
216 416
216 400
238 400
1 1 9 0 0 0 0 26 20 0 0 2
172 382
238 382
3 1 2 0 0 8320 0 37 31 0 0 2
440 276
487 276
3 1 3 0 0 4224 0 35 32 0 0 2
373 200
500 200
3 2 4 0 0 8320 0 34 37 0 0 3
372 299
372 285
394 285
3 1 5 0 0 12416 0 33 37 0 0 4
371 253
372 253
372 267
394 267
0 2 6 0 0 4096 0 0 33 43 0 2
296 262
326 262
0 1 7 0 0 4096 0 0 33 44 0 3
289 193
289 244
326 244
1 2 6 0 0 8320 0 28 35 0 0 4
173 324
296 324
296 209
324 209
3 1 7 0 0 20608 0 36 35 0 0 5
287 192
287 193
289 193
289 191
324 191
0 2 8 0 0 8192 0 0 34 47 0 3
191 217
191 308
327 308
0 1 9 0 0 4096 0 0 34 48 0 3
208 183
208 290
327 290
1 2 8 0 0 12416 0 29 36 0 0 4
174 217
216 217
216 201
238 201
1 1 9 0 0 4224 0 30 36 0 0 2
172 183
238 183
7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
438 646 489 667
447 653 479 668
4 Cout
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
434 451 485 472
443 458 475 473
4 Cout
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
433 252 484 273
442 259 474 274
4 Cout
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
449 375 484 396
458 382 474 397
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
454 570 489 591
463 577 479 592
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
456 771 489 792
464 778 480 793
2 S3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
439 175 474 196
448 182 464 197
2 S0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
