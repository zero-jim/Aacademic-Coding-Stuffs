CircuitMaker Text
5.6
Probes: 1
Q7_3
DC Sweep
0 339 244 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 130 30 200 10
1093 99 1909 1007
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
1261 195 2077 649
9961490 0
0
6 Title:
5 Name:
0
0
0
8
13 Logic Switch~
5 108 247 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8885 0 0
2
43535.1 2
0
14 Logic Display~
6 368 219 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3780 0 0
2
43535.1 7
0
2 +V
167 241 123 0 1 3
0 5
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9265 0 0
2
43535.1 6
0
7 Ground~
168 243 380 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9442 0 0
2
43535.1 5
0
9 N-MESFET~
219 288 305 0 3 7
0 6 3 2
0
0 0 848 0
7 NMESFET
11 0 60 8
2 Q8
29 -10 43 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
90 0 0 0 1 0 0 0
1 Q
9424 0 0
2
43535.1 4
0
9 P-MESFET~
219 288 184 0 3 7
0 5 3 6
0
0 0 848 0
7 PMESFET
11 0 60 8
2 Q7
29 -10 43 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
122 0 0 0 1 0 0 0
1 Q
9968 0 0
2
43535.1 3
0
9 P-MESFET~
219 183 186 0 3 7
0 5 4 3
0
0 0 848 0
7 PMESFET
11 0 60 8
2 Q4
29 -10 43 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
122 0 0 0 1 0 0 0
1 Q
9281 0 0
2
43535.1 1
0
9 N-MESFET~
219 183 307 0 3 7
0 3 4 2
0
0 0 848 0
7 NMESFET
11 0 60 8
2 Q3
29 -10 43 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
90 0 0 0 1 0 0 0
1 Q
8464 0 0
2
43535.1 0
0
11
0 0 3 0 0 4096 0 0 0 8 10 2
191 246
267 246
1 0 4 0 0 4112 0 1 0 0 7 2
120 247
162 247
1 0 5 0 0 4112 0 3 0 0 4 2
241 132
241 144
1 1 5 0 0 8336 0 6 7 0 0 4
296 166
296 144
191 144
191 168
3 0 2 0 0 8336 0 5 0 0 6 3
296 323
296 357
243 357
3 1 2 0 0 16 0 8 4 0 0 4
191 325
191 357
243 357
243 374
2 2 4 0 0 8336 0 7 8 0 0 4
170 186
162 186
162 307
170 307
3 1 3 0 0 4240 0 7 8 0 0 2
191 204
191 289
0 1 6 0 0 4112 0 0 2 11 0 3
296 245
368 245
368 237
2 2 3 0 0 8336 0 6 5 0 0 4
275 184
267 184
267 305
275 305
3 1 6 0 0 4240 0 6 5 0 0 2
296 202
296 287
0
0
2071 0 1
2 V4
0
2 V4
0 5 0.001
0
0 0 0
3 0 1 4
0 5e-06 2e-08 2e-08
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
