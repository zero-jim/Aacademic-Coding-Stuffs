CircuitMaker Text
5.6
Probes: 1
L1_1
DC Sweep
0 546 341 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
170 100 30 150 10
1093 99 1909 1007
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
1261 195 2077 649
9961490 0
0
6 Title:
5 Name:
0
0
0
11
13 Logic Switch~
5 231 379 0 1 11
0 6
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7876 0 0
2
43535.1 0
0
13 Logic Switch~
5 231 329 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6369 0 0
2
43535.1 1
0
9 P-MESFET~
219 504 280 0 3 7
0 5 4 3
0
0 0 848 0
7 PMESFET
11 0 60 8
2 Q6
29 -10 43 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
122 0 0 0 0 0 0 0
1 Q
9172 0 0
2
43535.1 0
0
9 N-MESFET~
219 504 401 0 3 7
0 3 4 2
0
0 0 848 0
7 NMESFET
11 0 60 8
2 Q5
29 -10 43 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
90 0 0 0 0 0 0 0
1 Q
7100 0 0
2
43535.1 0
0
7 Ground~
168 357 491 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3820 0 0
2
43535.1 2
0
2 +V
167 348 178 0 1 3
0 5
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7678 0 0
2
43535.1 3
0
14 Logic Display~
6 584 315 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
961 0 0
2
43535.1 4
0
9 N-MESFET~
219 433 425 0 3 7
0 4 7 2
0
0 0 848 512
7 NMESFET
-67 0 -18 8
2 Q4
-49 -10 -35 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
90 0 0 0 1 0 0 0
1 Q
3178 0 0
2
43535.1 5
0
9 N-MESFET~
219 289 426 0 3 7
0 4 6 2
0
0 0 848 0
7 NMESFET
11 0 60 8
2 Q3
29 -10 43 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
90 0 0 0 1 0 0 0
1 Q
3409 0 0
2
43535.1 6
0
9 P-MESFET~
219 340 274 0 3 7
0 8 7 4
0
0 0 848 0
7 PMESFET
11 0 60 8
2 Q2
29 -10 43 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
122 0 0 0 1 0 0 0
1 Q
3951 0 0
2
43535.1 7
0
9 P-MESFET~
219 340 223 0 3 7
0 5 6 8
0
0 0 848 0
7 PMESFET
11 0 60 8
2 Q1
29 -10 43 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
122 0 0 0 1 0 0 0
1 Q
8885 0 0
2
43535.1 8
0
16
0 1 3 0 0 4096 0 0 7 5 0 3
512 341
584 341
584 333
0 0 4 0 0 4224 0 0 0 3 11 2
483 341
348 341
2 2 4 0 0 0 0 3 4 0 0 4
491 280
483 280
483 401
491 401
3 0 2 0 0 8320 0 4 0 0 12 3
512 419
512 471
357 471
3 1 3 0 0 4240 0 3 4 0 0 2
512 298
512 383
1 0 5 0 0 8320 0 3 0 0 16 3
512 262
512 197
348 197
0 2 6 0 0 4224 0 0 11 10 0 3
272 379
272 223
327 223
0 2 7 0 0 4096 0 0 10 9 0 3
303 329
303 274
327 274
1 2 7 0 0 12416 0 2 8 0 0 6
243 329
303 329
303 378
449 378
449 425
440 425
1 2 6 0 0 0 0 1 9 0 0 4
243 379
273 379
273 426
276 426
0 3 4 0 0 0 0 0 10 14 0 2
348 399
348 292
1 0 2 0 0 0 0 5 0 0 13 2
357 485
357 451
3 3 2 0 0 128 0 9 8 0 0 4
297 444
297 451
419 451
419 443
1 1 4 0 0 128 0 9 8 0 0 4
297 408
297 399
419 399
419 407
1 3 8 0 0 4224 0 10 11 0 0 2
348 256
348 241
1 1 5 0 0 128 0 11 6 0 0 2
348 205
348 187
0
0
2071 0 1
2 V3
0
2 V3
0 5 0.001
0
0 0 0
3 0 1 4
0 5e-06 2e-08 2e-08
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
